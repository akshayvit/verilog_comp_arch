module andgate (x,y,z);
input x,y;
output z;
asign z=x&y;      
//similarly | for or gate and ~ for not 
endmodule